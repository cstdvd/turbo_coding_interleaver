configuration cfg of interleaver_tb is
	for interleaver_test
		-- configurazione di default
	end for;
end cfg;
